module adder (
    input  data_1_i,
    input  data_2_i,
    output sum_o
);
    assign sum_o = data_1_i + data_2_i;
endmodule
